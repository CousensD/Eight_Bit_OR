module tt_um_or(
  input clk,
  input reset,
  input [7:0] a, b,
  output [7:0] Y
);

  assign Y = a | b;

  endmodule
    
